module InstBuffer (
    
);
    
endmodule